module carry_select_adder ();

endmodule
