// add/sub/div/divu/mul/mulu
// clo (leading ones)
// clz (leading zeros)
// low2high
// low2low
// hight2low
//
module alu ();

endmodule
