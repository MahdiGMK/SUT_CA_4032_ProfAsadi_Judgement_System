module carry_select_adder #(
    parameter int N = 32
) (
    input [N-1:0] a,
    input [N-1:0] b,
    input cin,
    output [N-1:0] s,
    output cout
);

endmodule
